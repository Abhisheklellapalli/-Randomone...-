class transaction;
  randc bit rst;
  randc bit t;
endclass
