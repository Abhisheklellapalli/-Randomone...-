interface dff;
  logic clk,rst;
  logic d;
  logic q;
  logic qbar;
endinterface
