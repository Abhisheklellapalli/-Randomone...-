class trans;
  rand bit j;
  rand bit k;
  rand bit rst;
endclass
