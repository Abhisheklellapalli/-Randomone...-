class transaction;
  rand bit d;
  randc bit rst;
endclass
