interface ff;
  reg clk;
  reg rst;
  reg t;
  reg q;
  reg qbar;
endinterface
