typedef struct{ 
  bit a;     //demux input
  logic [1:0] s; //selection lines
  logic [3:0]y; // output
} value_s;
