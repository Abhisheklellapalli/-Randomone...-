// _____________________________________
// |                                   |
// |          RANDOM K MAP             |
// |___________________________________|
//      00     01      11      10    
//   --------------------------------
//   |      |       |       |       |
// 0 |      |   1   |       |  1    |
//   |      |       |       |       |
//   -------+-------+-------+--------
//   |      |       |       |       |
// 1 |  1   |   1   |   1   |       |
//   |      |       |       |       |
//   --------------------------------
// F(A,B,C) = A(B'+C)+A'BC'+B'C

module kmap(
  input a,b,c,
  output f
);
  assign f = (a&(~b|c))|(~a&b&~c)|~b&c;
endmodule
