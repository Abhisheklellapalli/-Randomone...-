interface dm;
  logic a;
  logic [1:0]s;
  logic [3:0]y;
endinterface
