typedef struct { 
  bit a,b,borin;
  bit dif,borout;
} ports;
