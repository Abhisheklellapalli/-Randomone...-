module encoder_32_to_5_tb;
    reg [31:0] in;
    wire [4:0] out;
 encoder_32_to_5 haa( .in(in), .out(out));
 initial
 begin
$display("Time\t\tInput Bit\tOutput");
$monitor("%0t\t%b\t%0d", $time, in, out);
   
   in =32'b00000000000000000000000000000001;
   #10;
   in =32'b00000000000000000000000000000010;
   #10;
   in =32'b00000000000000000000000000000100;
   #10;
   in =32'b00000000000000000000000000001000;
   #10;
   in =32'b00000000000000000000000000010000;
   #10;
   in =32'b00000000000000000000000000100000;
   #10;
   in =32'b00000000000000000000000001000000;
   #10;
   in =32'b00000000000000000000000010000000;
   #10;
   in =32'b00000000000000000000000100000000;
   #10;
   in =32'b00000000000000000000001000000000;
   #10;
   in =32'b00000000000000000000010000000000;
   #10;
   in =32'b00000000000000000000100000000000;
   #10;
   in =32'b00000000000000000001000000000000;
   #10;
   in =32'b00000000000000000010000000000000;
   #10;
   in =32'b00000000000000000100000000000000;
   #10;
   in =32'b00000000000000001000000000000000;
   #10;
   in =32'b00000000000000010000000000000000;
   #10;
   in =32'b00000000000000100000000000000000;
   #10;
   in =32'b00000000000001000000000000000000;
   #10;
   in =32'b00000000000010000000000000000000;
   #10;
   in =32'b00000000000100000000000000000000;
   #10;
   in =32'b00000000001000000000000000000000;
   #10;
   in =32'b00000000010000000000000000000000;
   #10;
   in =32'b00000000100000000000000000000000;
   #10;
   in =32'b00000001000000000000000000000000;
   #10;
   in =32'b00000010000000000000000000000000;
   #10;
   in =32'b00000100000000000000000000000000;
   #10;
   in =32'b00001000000000000000000000000000;
   #10;
   in =32'b00010000000000000000000000000000;
   #10;
   in =32'b00100000000000000000000000000000;
   #10;
   in =32'b01000000000000000000000000000000;
   #10;
   in =32'b10000000000000000000000000000000;
   #10;
 $finish;
 
 end
endmodule
