// Interface
interface fs;
  logic a,b,borin;
  logic dif,borout;
endinterface
