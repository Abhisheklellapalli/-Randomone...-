class transaction;
  randc bit rst;
  rand bit s;
  rand bit r;
endclass
