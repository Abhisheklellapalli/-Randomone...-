// interface 

interface hs;
  logic a,b;
  logic diff,bor;
endinterface
