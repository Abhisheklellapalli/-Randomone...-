interface srff;
  logic clk;
  logic rst;
  logic s;
  logic r;
  logic q;
  logic qbar;
endinterface
