interface j_k_ff;
  logic clk;
  logic rst;
  logic j;
  logic k;
  logic q;
  logic qbar;
endinterface
